library verilog;
use verilog.vl_types.all;
entity socket_txd is
    generic(
        IDLE            : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        RDFSR_CMD       : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        RD_FSR          : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        JDFSR           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        WRIR_CMD        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        WR_IR           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        RDTXWD_CMD      : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        RD_TX_WD        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        WRDIP_CMD       : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        WR_DIP          : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        WRDPORT_CMD     : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        WR_DPORT        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        WRTXBUF_CMD     : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi0);
        WR_TXBUF        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi1);
        WRTXWD_CMD      : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        WR_TXWD         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        WRCR_CMD        : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        WR_CR           : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        RDIR_CMD        : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi0);
        RD_IR           : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi1);
        JDIR            : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi0);
        \END\           : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi1);
        SN_DIP          : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        SN_DPORT        : vl_logic_vector(0 to 15) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        SN_DSHAR        : vl_logic_vector(0 to 47) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        SN_PORT         : vl_logic_vector(0 to 15) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        rdreq           : in     vl_logic;
        den             : in     vl_logic;
        din             : in     vl_logic_vector(7 downto 0);
        task_state      : in     vl_logic_vector(3 downto 0);
        txdat_vld       : in     vl_logic;
        txdat           : in     vl_logic_vector(7 downto 0);
        txdat_len       : in     vl_logic_vector(15 downto 0);
        dat_tx_req      : in     vl_logic;
        o_dat_rx_rden   : out    vl_logic;
        wrend           : in     vl_logic;
        o_start         : out    vl_logic;
        o_cmd           : out    vl_logic_vector(7 downto 0);
        o_addr          : out    vl_logic_vector(15 downto 0);
        o_length        : out    vl_logic_vector(15 downto 0);
        o_dat           : out    vl_logic_vector(7 downto 0);
        o_tx_end        : out    vl_logic;
        o_ts            : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of RDFSR_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_FSR : constant is 1;
    attribute mti_svvh_generic_type of JDFSR : constant is 1;
    attribute mti_svvh_generic_type of WRIR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_IR : constant is 1;
    attribute mti_svvh_generic_type of RDTXWD_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_TX_WD : constant is 1;
    attribute mti_svvh_generic_type of WRDIP_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_DIP : constant is 1;
    attribute mti_svvh_generic_type of WRDPORT_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_DPORT : constant is 1;
    attribute mti_svvh_generic_type of WRTXBUF_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_TXBUF : constant is 1;
    attribute mti_svvh_generic_type of WRTXWD_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_TXWD : constant is 1;
    attribute mti_svvh_generic_type of WRCR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_CR : constant is 1;
    attribute mti_svvh_generic_type of RDIR_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_IR : constant is 1;
    attribute mti_svvh_generic_type of JDIR : constant is 1;
    attribute mti_svvh_generic_type of \END\ : constant is 1;
    attribute mti_svvh_generic_type of SN_DIP : constant is 1;
    attribute mti_svvh_generic_type of SN_DPORT : constant is 1;
    attribute mti_svvh_generic_type of SN_DSHAR : constant is 1;
    attribute mti_svvh_generic_type of SN_PORT : constant is 1;
end socket_txd;

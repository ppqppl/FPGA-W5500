library verilog;
use verilog.vl_types.all;
entity ini_w5500 is
    generic(
        GAR             : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        SUBR            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SHAR            : vl_logic_vector(0 to 47) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        SIPR            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        IDLE            : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RST             : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        WRMR_CMD        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        WR_MR           : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        RDMR_CMD        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        RD_MR           : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        JDMR            : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        WRGAR_CMD       : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        WR_GAR          : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        WRSUBR_CMD      : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        WR_SUBR         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        WRSHAR_CMD      : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        WR_SHAR         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        WRIP_CMD        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        WR_IP           : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        RDRG_CMD        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        RD_RG           : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        JDRG            : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        WRIR_CMD        : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        WR_IR           : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        WRIMR_CMD       : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        WR_IMR          : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        RDIR_CMD        : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        RD_IR           : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        JDIR            : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        WRRTR_CMD       : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        WR_RTR          : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        RDRTR_CMD       : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        RD_RTR          : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        JDRTR           : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        WRRCR_CMD       : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        WR_RCR          : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        RDRCR_CMD       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        RD_RCR          : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        JDRCR           : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        WRPHY_CMD       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        WR_PHY          : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        RDPHY_CMD       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        RD_PHY          : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        JDPHY           : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        \END\           : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        RSTNUM          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        DLYNUM          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0)
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        ini_en          : in     vl_logic;
        rdreq           : in     vl_logic;
        den             : in     vl_logic;
        din             : in     vl_logic_vector(7 downto 0);
        wrend           : in     vl_logic;
        o_start         : out    vl_logic;
        o_cmd           : out    vl_logic_vector(7 downto 0);
        o_addr          : out    vl_logic_vector(15 downto 0);
        o_length        : out    vl_logic_vector(15 downto 0);
        o_dat           : out    vl_logic_vector(7 downto 0);
        o_w5500_rst     : out    vl_logic;
        o_ini_end       : out    vl_logic;
        o_ts            : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GAR : constant is 1;
    attribute mti_svvh_generic_type of SUBR : constant is 1;
    attribute mti_svvh_generic_type of SHAR : constant is 1;
    attribute mti_svvh_generic_type of SIPR : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of RST : constant is 1;
    attribute mti_svvh_generic_type of WRMR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_MR : constant is 1;
    attribute mti_svvh_generic_type of RDMR_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_MR : constant is 1;
    attribute mti_svvh_generic_type of JDMR : constant is 1;
    attribute mti_svvh_generic_type of WRGAR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_GAR : constant is 1;
    attribute mti_svvh_generic_type of WRSUBR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_SUBR : constant is 1;
    attribute mti_svvh_generic_type of WRSHAR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_SHAR : constant is 1;
    attribute mti_svvh_generic_type of WRIP_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_IP : constant is 1;
    attribute mti_svvh_generic_type of RDRG_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_RG : constant is 1;
    attribute mti_svvh_generic_type of JDRG : constant is 1;
    attribute mti_svvh_generic_type of WRIR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_IR : constant is 1;
    attribute mti_svvh_generic_type of WRIMR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_IMR : constant is 1;
    attribute mti_svvh_generic_type of RDIR_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_IR : constant is 1;
    attribute mti_svvh_generic_type of JDIR : constant is 1;
    attribute mti_svvh_generic_type of WRRTR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_RTR : constant is 1;
    attribute mti_svvh_generic_type of RDRTR_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_RTR : constant is 1;
    attribute mti_svvh_generic_type of JDRTR : constant is 1;
    attribute mti_svvh_generic_type of WRRCR_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_RCR : constant is 1;
    attribute mti_svvh_generic_type of RDRCR_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_RCR : constant is 1;
    attribute mti_svvh_generic_type of JDRCR : constant is 1;
    attribute mti_svvh_generic_type of WRPHY_CMD : constant is 1;
    attribute mti_svvh_generic_type of WR_PHY : constant is 1;
    attribute mti_svvh_generic_type of RDPHY_CMD : constant is 1;
    attribute mti_svvh_generic_type of RD_PHY : constant is 1;
    attribute mti_svvh_generic_type of JDPHY : constant is 1;
    attribute mti_svvh_generic_type of \END\ : constant is 1;
    attribute mti_svvh_generic_type of RSTNUM : constant is 1;
    attribute mti_svvh_generic_type of DLYNUM : constant is 1;
end ini_w5500;

library verilog;
use verilog.vl_types.all;
entity ama_systolic_adder_function is
    generic(
        width_data_in   : integer := 1;
        width_chainin   : integer := 1;
        width_data_out  : integer := 1;
        number_of_adder_input: integer := 1;
        systolic_delay1 : string  := "UNREGISTERED";
        systolic_aclr1  : string  := "NONE";
        systolic_delay3 : string  := "UNREGISTERED";
        systolic_aclr3  : string  := "NONE";
        adder1_direction: string  := "NONE";
        adder3_direction: string  := "NONE";
        port_addnsub1   : string  := "PORT_UNUSED";
        addnsub_multiplier_register1: string  := "CLOCK0";
        addnsub_multiplier_aclr1: string  := "ACLR3";
        port_addnsub3   : string  := "PORT_UNUSED";
        addnsub_multiplier_register3: string  := "CLOCK0";
        addnsub_multiplier_aclr3: string  := "ACLR3";
        latency         : integer := 0;
        addnsub_multiplier_latency_clock1: string  := "UNREGISTERED";
        addnsub_multiplier_latency_aclr1: string  := "NONE";
        addnsub_multiplier_latency_clock3: string  := "UNREGISTERED";
        addnsub_multiplier_latency_aclr3: string  := "NONE";
        width_data_in_msb: vl_notype;
        width_data_out_msb: vl_notype;
        width_chainin_msb: vl_notype;
        width_systolic  : vl_notype;
        width_systolic_msb: vl_notype;
        input_ext_width : vl_notype
    );
    port(
        data_in_0       : in     vl_logic_vector;
        data_in_1       : in     vl_logic_vector;
        data_in_2       : in     vl_logic_vector;
        data_in_3       : in     vl_logic_vector;
        chainin         : in     vl_logic_vector;
        clock           : in     vl_logic_vector(3 downto 0);
        aclr            : in     vl_logic_vector(3 downto 0);
        ena             : in     vl_logic_vector(3 downto 0);
        data_out        : out    vl_logic_vector;
        addnsub1        : in     vl_logic;
        addnsub3        : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width_data_in : constant is 1;
    attribute mti_svvh_generic_type of width_chainin : constant is 1;
    attribute mti_svvh_generic_type of width_data_out : constant is 1;
    attribute mti_svvh_generic_type of number_of_adder_input : constant is 1;
    attribute mti_svvh_generic_type of systolic_delay1 : constant is 1;
    attribute mti_svvh_generic_type of systolic_aclr1 : constant is 1;
    attribute mti_svvh_generic_type of systolic_delay3 : constant is 1;
    attribute mti_svvh_generic_type of systolic_aclr3 : constant is 1;
    attribute mti_svvh_generic_type of adder1_direction : constant is 1;
    attribute mti_svvh_generic_type of adder3_direction : constant is 1;
    attribute mti_svvh_generic_type of port_addnsub1 : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_register1 : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_aclr1 : constant is 1;
    attribute mti_svvh_generic_type of port_addnsub3 : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_register3 : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_aclr3 : constant is 1;
    attribute mti_svvh_generic_type of latency : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_latency_clock1 : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_latency_aclr1 : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_latency_clock3 : constant is 1;
    attribute mti_svvh_generic_type of addnsub_multiplier_latency_aclr3 : constant is 1;
    attribute mti_svvh_generic_type of width_data_in_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_out_msb : constant is 3;
    attribute mti_svvh_generic_type of width_chainin_msb : constant is 3;
    attribute mti_svvh_generic_type of width_systolic : constant is 3;
    attribute mti_svvh_generic_type of width_systolic_msb : constant is 3;
    attribute mti_svvh_generic_type of input_ext_width : constant is 3;
end ama_systolic_adder_function;
